library ieee;
use ieee.std_logic_1164.all;
entity coeffs is
port( b : out std_logic_vector(383 downto 0));
end entity;
architecture behavioral of coeffs is
begin
"000000000101",
"000000000110",
"000000001001",
"000000001110",
"000000010101",
"000000011101",
"000000101000",
"000000110100",
"000001000001",
"000001001111",
"000001011100",
"000001101001",
"000001110100",
"000001111101",
"000010000011",
"000010000110",
"000010000110",
"000010000011",
"000001111101",
"000001110100",
"000001101001",
"000001011100",
"000001001111",
"000001000001",
"000000110100",
"000000101000",
"000000011101",
"000000010101",
"000000001110",
"000000001001",
"000000000110",
"000000000101",
end architecture behavioral;
